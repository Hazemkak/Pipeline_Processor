Library ieee;
use ieee.std_logic_1164.all;

entity control is 
PORT
( op_code: IN std_logic_vector(4 DOWNTO 0);
control_signals : OUT std_logic_vector(25 DOWNTO 0)
);
END control;

architecture archcontrol of control is
    begin
  
    with op_code select
    control_signals <= 
            "00000000000000001000000000" when "00000",
            "00000000000000001000000000" when "00001",
            "00000000000000001000100010" when "00010",
            "00001000000000001001000101" when "00011",
            "00001000000000001001100111" when "00100",
            "00000010000000001000000001" when "00101",
            "00001100000000001000000000" when "00110",
            "00001000000000001000000001" when "00111",
            "00001000000000001001101001" when "01000",
            "00001000000000001001101011" when "01001",
            "00001000000000001001001101" when "01010",
            "00001000000000001001111001" when "01011",
            "00100000000100001000000001" when "01100",
            "01111000001000001000000000" when "01101",
            "00001000000000001000010000" when "01110",
            "00011000001000001000011001" when "01111",
            "00000000000100001000011001" when "10000",
            "00000000000000001000000000" when others;
            
   
  
end archcontrol ;